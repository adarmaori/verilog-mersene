module divisibility_checker (
  input clk,
  input a,
  input b,
  output done,
  output divisible
);
  
endmodule
